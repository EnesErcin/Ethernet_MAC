module transmit_controller (
    
    input gmii_buffer_full,
    output logic gmii_tx_en
    output logic gmii_clk,
);
    
endmodule