package global;
  parameter initial_value = 1;
  parameter crc_len = 32;
  parameter crc_poly = 32'h04C11DB7;
  parameter datalen = 8;
  parameter payload_len = 11'd9;
endpackage