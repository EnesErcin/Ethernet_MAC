
package utils;
    parameter  min_payload_len =                 16'd46;
    parameter  len_addr        =                 13'd6;
    parameter  len_len         =                 13'd2;
    parameter  len_crc         =                 13'd4;
    parameter  len_perm        =                 13'd7;
    parameter  len_max_payload =                 50;
endpackage

