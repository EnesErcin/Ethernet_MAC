`define min_payload_len 16'd46
`define len_addr    13'd6
`define len_len     13'd2
`define len_crc     13'd4
`define len_perm    13'd7